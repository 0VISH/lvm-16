module not16(output wire [15:0] out, input wire [15:0] in);

assign out = ~in;

endmodule;
